module xor_gate(input q,t, output y  );

assign y= q ^ t;

endmodule