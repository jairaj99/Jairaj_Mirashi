package ahb_apb_pkg;

    import uvm_pkg::*;
        
		`include "uvm_macros.svh"
		
        `include "ahb_config.sv"
        `include "ahb_driver.sv"
        `include "ahb_monitor.sv"
        `include "ahb_agent.sv"
        `include "ahb_agt_top.sv"

		`include "apb_config.sv"
        `include "apb_driver.sv"
        `include "apb_monitor.sv"
        `include "apb_agent.sv"
        `include "apb_agt_top.sv"
		
		`include "ahb_apb_env_config.sv"
        `include "ahb_apb_env.sv"


endpackage