// Define the interface not_if
interface not_if();
  // Declare the signals in the interface
  logic in;  // Input signal for the DUT
  logic out; // Output signal from the DUT
endinterface
